module encoder8_3_tb;
  reg [7:0] d;
  wire [2:0] y;
  encoder8_3 en(d,y);
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(1);
    d[0]=1;d[1]=0;d[2]=0;d[3]=0;d[4]=0;d[5]=0;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=1;d[2]=0;d[3]=0;d[4]=0;d[5]=0;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=1;d[3]=0;d[4]=0;d[5]=0;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=0;d[3]=1;d[4]=0;d[5]=0;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=0;d[3]=0;d[4]=1;d[5]=0;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=0;d[3]=0;d[4]=0;d[5]=1;d[6]=0;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=0;d[3]=0;d[4]=0;d[5]=0;d[6]=1;d[7]=0;#5
    d[0]=0;d[1]=0;d[2]=0;d[3]=0;d[4]=0;d[5]=0;d[6]=0;d[7]=1;#5

    $finish;
 
  
  end
endmodule
